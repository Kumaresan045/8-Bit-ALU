module NOT(input [7:0] op1, output [7:0] res); //8-bit bitwise NOT

    not modulei[7:0] (res[7:0], op1[7:0]);

endmodule
